/*
Author: Sajeed Mohammad Shahriat
Affiliation: Rochester Institute of Technology
All rights reserved
This files can be reused and modified given that this copyright notice is not removed
*/

module hello_world;

initial
	begin
		$display ("Hello World");
		#10
		$finish;
	end
endmodule
